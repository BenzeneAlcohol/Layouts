*nmos inverter with resistive load

.include ./t14y_tsmc_025_level3.txt

*netlist
m0 x in 0 0 cmosn w=2u l=1u
rl vdd out 10k
cl y 0 1f

*voltage sources
v_dd vdd 0 dc 5
v_x out x dc 0
v_in in 0 dc 5 pulse(0 5 1n 0.1n 0.1n 2n 4n)
v_y out y dc 0

*analysis
.control
	foreach wid 5u 10u 20u
		alter m0 w=$wid
		
		dc v_in 0 5 0.1
		setplot dc$wid
		plot in out
		
		tran 0.1n 6n
		meas tran vmin MIN out from=1.9n to=2.1n
		meas tran vmax MAX out from=3.9n to=4.1n
		
		let v10 = vmin + 0.1*(vmax - vmin)
		let v50 = vmin + 0.5*(vmax - vmin)
		let v90 = vmin + 0.9*(vmax - vmin)
		
		meas tran trise trig out val=v10 rise=1 targ out val=v90 rise=1
		meas tran tfall trig out val=v90 fall=1 targ out val=v10 fall=1
		
		meas tran tplh trig in val=2.5 fall=1 targ out val=v50 rise=1
		meas tran tphl trig in val=2.5 rise=1 targ out val=v50 fall=1
		
		let tp = 0.5*(tplh + tphl)

		let power = vdd * (-v_x#branch)
		meas tran avg_pow AVG power from=2n to=6n	
				
		print vmin vmax trise tfall tp avg_pow
	end
		
.endc

.end
