magic
tech scmos
timestamp 1667411863
<< nwell >>
rect -19 21 8 47
<< polysilicon >>
rect -13 32 -11 34
rect 0 32 2 34
rect -13 18 -11 22
rect -20 14 -11 18
rect -13 9 -11 14
rect 0 18 2 22
rect 0 14 10 18
rect 0 9 2 14
rect -13 -3 -11 -1
rect 0 -3 2 -1
<< ndiffusion >>
rect -14 5 -13 9
rect -18 -1 -13 5
rect -11 -1 0 9
rect 2 5 3 9
rect 2 -1 7 5
<< pdiffusion >>
rect -14 28 -13 32
rect -18 22 -13 28
rect -11 26 0 32
rect -11 22 -8 26
rect -4 22 0 26
rect 2 28 3 32
rect 2 22 7 28
<< metal1 >>
rect -18 45 7 46
rect -18 41 -7 45
rect -3 41 7 45
rect -18 40 7 41
rect -18 32 -14 40
rect 3 32 7 40
rect -8 18 -4 22
rect -8 13 7 18
rect 3 9 7 13
rect -18 -9 -14 5
rect -18 -10 7 -9
rect -18 -14 -8 -10
rect -4 -14 7 -10
rect -18 -15 7 -14
<< ntransistor >>
rect -13 -1 -11 9
rect 0 -1 2 9
<< ptransistor >>
rect -13 22 -11 32
rect 0 22 2 32
<< polycontact >>
rect -24 14 -20 18
rect 10 14 14 18
<< ndcontact >>
rect -18 5 -14 9
rect 3 5 7 9
<< pdcontact >>
rect -18 28 -14 32
rect -8 22 -4 26
rect 3 28 7 32
<< psubstratepcontact >>
rect -8 -14 -4 -10
<< nsubstratencontact >>
rect -7 41 -3 45
<< labels >>
rlabel metal1 3 41 7 45 3 vdd
rlabel metal1 3 -14 7 -10 3 vss
rlabel polycontact 10 14 14 18 3 vin_b
rlabel polycontact -24 14 -20 18 7 vin_a
rlabel metal1 -8 14 -4 18 5 vout
<< end >>
