magic
tech scmos
timestamp 1667332312
<< nwell >>
rect -5 -33 14 2
<< polysilicon >>
rect 2 -12 7 -10
rect 2 -37 7 -32
rect -5 -41 7 -37
rect 2 -46 7 -41
rect 2 -58 7 -56
<< ndiffusion >>
rect 0 -50 2 -46
rect -4 -56 2 -50
rect 7 -50 9 -46
rect 7 -56 13 -50
<< pdiffusion >>
rect -4 -28 2 -12
rect 0 -32 2 -28
rect 7 -28 13 -12
rect 7 -32 9 -28
<< metal1 >>
rect -4 -3 8 1
rect 12 -3 13 1
rect -4 -4 13 -3
rect -4 -28 0 -4
rect 9 -46 13 -32
rect -4 -65 0 -50
rect -4 -69 8 -65
rect 12 -69 13 -65
rect -4 -70 13 -69
<< ntransistor >>
rect 2 -56 7 -46
<< ptransistor >>
rect 2 -32 7 -12
<< polycontact >>
rect -9 -41 -5 -37
<< ndcontact >>
rect -4 -50 0 -46
rect 9 -50 13 -46
<< pdcontact >>
rect -4 -32 0 -28
rect 9 -32 13 -28
<< psubstratepcontact >>
rect 8 -69 12 -65
<< nsubstratencontact >>
rect 8 -3 12 1
<< labels >>
rlabel polycontact -9 -41 -5 -37 7 vin
rlabel metal1 9 -41 13 -37 3 vout
rlabel metal1 1 -3 5 1 1 vdd
rlabel metal1 1 -70 5 -66 5 vss
<< end >>
