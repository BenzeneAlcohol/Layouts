magic
tech scmos
timestamp 1667423039
<< nwell >>
rect -11 1 31 21
<< polysilicon >>
rect -4 12 -2 14
rect 12 12 14 14
rect 22 12 24 14
rect -4 0 -2 2
rect -9 -4 -2 0
rect -4 -14 -2 -4
rect 12 -1 14 2
rect 12 -5 15 -1
rect 12 -14 14 -5
rect 22 -7 24 2
rect 22 -11 33 -7
rect 22 -14 24 -11
rect -4 -26 -2 -24
rect 12 -26 14 -24
rect 22 -26 24 -24
<< ndiffusion >>
rect -10 -20 -4 -14
rect -6 -24 -4 -20
rect -2 -24 12 -14
rect 14 -24 22 -14
rect 24 -18 26 -14
rect 24 -24 30 -18
<< pdiffusion >>
rect -6 8 -4 12
rect -10 2 -4 8
rect -2 6 12 12
rect -2 2 0 6
rect 4 2 12 6
rect 14 8 16 12
rect 20 8 22 12
rect 14 2 22 8
rect 24 6 30 12
rect 24 2 26 6
<< metal1 >>
rect -10 16 0 20
rect 4 16 20 20
rect -10 12 -6 16
rect 16 12 20 16
rect 0 -8 4 2
rect 26 -8 30 2
rect 0 -12 30 -8
rect 26 -14 30 -12
rect -10 -30 -6 -24
rect -10 -31 24 -30
rect -10 -35 2 -31
rect 6 -35 24 -31
<< ntransistor >>
rect -4 -24 -2 -14
rect 12 -24 14 -14
rect 22 -24 24 -14
<< ptransistor >>
rect -4 2 -2 12
rect 12 2 14 12
rect 22 2 24 12
<< polycontact >>
rect -13 -4 -9 0
rect 15 -5 19 -1
rect 33 -11 37 -7
<< ndcontact >>
rect -10 -24 -6 -20
rect 26 -18 30 -14
<< pdcontact >>
rect -10 8 -6 12
rect 0 2 4 6
rect 16 8 20 12
rect 26 2 30 6
<< psubstratepcontact >>
rect 2 -35 6 -31
<< nsubstratencontact >>
rect 0 16 4 20
<< labels >>
rlabel polycontact -13 -4 -9 0 7 vin_a
rlabel metal1 14 16 18 20 1 vdd
rlabel metal1 13 -35 17 -31 5 vss
rlabel polycontact 33 -11 37 -7 3 vin_c
rlabel polycontact 15 -5 19 -1 1 vin_b
rlabel metal1 26 -5 30 -1 3 vout
<< end >>
