magic
tech scmos
timestamp 1667372487
<< nwell >>
rect -8 7 14 60
<< polysilicon >>
rect -2 48 0 50
rect 6 48 8 50
rect -2 4 0 8
rect -8 0 0 4
rect -2 -4 0 0
rect 6 4 8 8
rect 6 0 16 4
rect 6 -4 8 0
rect -2 -16 0 -14
rect 6 -16 8 -14
<< ndiffusion >>
rect -7 -10 -2 -4
rect -3 -14 -2 -10
rect 0 -8 1 -4
rect 5 -8 6 -4
rect 0 -14 6 -8
rect 8 -10 13 -4
rect 8 -14 9 -10
<< pdiffusion >>
rect -3 44 -2 48
rect -7 8 -2 44
rect 0 8 6 48
rect 8 12 13 48
rect 8 8 9 12
<< metal1 >>
rect -7 58 13 59
rect -7 54 8 58
rect 12 54 13 58
rect -7 53 13 54
rect -7 48 -3 53
rect 9 4 13 8
rect 1 0 13 4
rect 1 -4 5 0
rect -7 -19 -3 -14
rect 9 -19 13 -14
rect -7 -25 13 -19
<< ntransistor >>
rect -2 -14 0 -4
rect 6 -14 8 -4
<< ptransistor >>
rect -2 8 0 48
rect 6 8 8 48
<< polycontact >>
rect -12 0 -8 4
rect 16 0 20 4
<< ndcontact >>
rect -7 -14 -3 -10
rect 1 -8 5 -4
rect 9 -14 13 -10
<< pdcontact >>
rect -7 44 -3 48
rect 9 8 13 12
<< nsubstratencontact >>
rect 8 54 12 58
<< labels >>
rlabel metal1 1 -24 5 -20 5 vss
rlabel metal1 1 0 5 4 1 vout
rlabel polycontact -12 0 -8 4 7 vin_a
rlabel polycontact 16 0 20 4 3 vin_b
rlabel metal1 1 54 5 58 1 vdd
<< end >>
