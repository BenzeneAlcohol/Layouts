* SPICE3 file created from func.ext - technology: scmos

.option scale=1u

M1000 vout vin_c a_n8_15# vdd pfet w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1001 vout vin_b a_0_n13# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 a_n8_15# vin_b vdd vdd pfet w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_0_n13# vin_a vss Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 vdd vin_a a_n8_15# vdd pfet w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 vss vin_c vout Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vss 0 7.52fF **FLOATING
C1 vout 0 4.70fF **FLOATING
C2 a_n8_15# 0 4.14fF **FLOATING
C3 vin_c 0 10.53fF **FLOATING
C4 vin_b 0 7.06fF **FLOATING
C5 vin_a 0 8.95fF **FLOATING
