magic
tech scmos
timestamp 1667421450
<< nwell >>
rect -13 12 26 38
<< polysilicon >>
rect -7 23 -5 25
rect 3 23 5 25
rect 14 23 16 25
rect -7 7 -5 13
rect -22 3 -5 7
rect -7 -8 -5 3
rect 3 5 5 13
rect 3 1 6 5
rect 3 -8 5 1
rect 14 -8 16 13
rect 21 4 25 8
rect -7 -20 -5 -18
rect 3 -20 5 -18
rect 14 -20 16 -18
<< ndiffusion >>
rect -12 -14 -7 -8
rect -8 -18 -7 -14
rect -5 -18 3 -8
rect 5 -18 14 -8
rect 16 -12 17 -8
rect 21 -12 25 -8
rect 16 -18 25 -12
<< pdiffusion >>
rect -8 19 -7 23
rect -12 13 -7 19
rect -5 17 3 23
rect -5 13 -3 17
rect 1 13 3 17
rect 5 19 8 23
rect 12 19 14 23
rect 5 13 14 19
rect 16 17 25 23
rect 16 13 17 17
rect 21 13 25 17
<< metal1 >>
rect -12 33 17 37
rect 21 33 25 37
rect -12 29 25 33
rect -12 23 -8 29
rect 8 23 12 29
rect -3 -2 1 13
rect 17 -2 21 13
rect -3 -6 21 -2
rect 17 -8 21 -6
rect -12 -25 -8 -18
rect -12 -26 25 -25
rect -12 -30 16 -26
rect 20 -30 25 -26
rect -12 -33 25 -30
<< ntransistor >>
rect -7 -18 -5 -8
rect 3 -18 5 -8
rect 14 -18 16 -8
<< ptransistor >>
rect -7 13 -5 23
rect 3 13 5 23
rect 14 13 16 23
<< polycontact >>
rect -26 3 -22 7
rect 6 1 10 5
rect 25 4 29 8
<< ndcontact >>
rect -12 -18 -8 -14
rect 17 -12 21 -8
<< pdcontact >>
rect -12 19 -8 23
rect -3 13 1 17
rect 8 19 12 23
rect 17 13 21 17
<< psubstratepcontact >>
rect 16 -30 20 -26
<< nsubstratencontact >>
rect 17 33 21 37
<< labels >>
rlabel metal1 2 33 6 37 1 vdd
rlabel polycontact 6 1 10 5 3 vin_b
rlabel polycontact 25 4 29 8 3 vin_c
rlabel metal1 4 -32 8 -28 5 vss
rlabel metal1 -3 -6 1 -2 7 vout
rlabel polycontact -26 3 -22 7 7 vin_a
<< end >>
