*nmos varying threshold voltage

.include t14y_tsmc_025_level3.txt

*netlist
m0 vdd in vss vss cmosn l=1u w=2u

*voltage sources declaration
v_dd vdd 0 dc 5
v_ss vss 0 dc 0
v_in in 0 dc 5

*analysis
.control
	foreach vth 0.2 1.0 1.5
		altermod m0 VTO = $vth
		
		dc v_in 0 5 0.1
		
		setplot dc$vth
		plot -v_dd#branch
		
	end
.endc

.end
	
	
