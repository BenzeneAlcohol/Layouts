*nmos characteristics varying vsb

.include ./t14y_tsmc_025_level3.txt

*netlist
m0 vdd in vss vbb cmosn l=1u w=2u

*voltage sources
v_dd vdd 0 dc 5
v_in in 0 dc 5
v_ss vss 0 dc 0
v_sb vss vbb dc 3


*analysis
.control
	dc v_in 0 5 0.1 v_sb 0 3 1
	
	setplot dc1
	plot -v_dd#branch
.endc

.end	





