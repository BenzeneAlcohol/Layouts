magic
tech scmos
timestamp 1667423900
<< nwell >>
rect -12 7 25 39
<< polysilicon >>
rect -5 28 -3 30
rect 5 28 7 30
rect 15 28 17 30
rect -5 2 -3 8
rect 5 5 7 8
rect -15 -2 -3 2
rect 4 1 7 5
rect -5 -10 -3 -2
rect 5 -10 7 1
rect 15 2 17 8
rect 15 -2 24 2
rect 15 -10 17 -2
rect -5 -22 -3 -20
rect 5 -22 7 -20
rect 15 -22 17 -20
<< ndiffusion >>
rect -7 -14 -5 -10
rect -11 -20 -5 -14
rect -3 -16 5 -10
rect -3 -20 -1 -16
rect 3 -20 5 -16
rect 7 -14 9 -10
rect 13 -14 15 -10
rect 7 -20 15 -14
rect 17 -16 24 -10
rect 17 -20 19 -16
rect 23 -20 24 -16
<< pdiffusion >>
rect -11 12 -5 28
rect -7 8 -5 12
rect -3 8 5 28
rect 7 8 15 28
rect 17 24 19 28
rect 23 24 24 28
rect 17 8 24 24
<< metal1 >>
rect -11 34 3 38
rect 7 34 23 38
rect -11 33 23 34
rect 19 28 23 33
rect -11 -4 -7 8
rect -11 -8 13 -4
rect -11 -10 -7 -8
rect 9 -10 13 -8
rect -1 -24 3 -20
rect 19 -24 23 -20
rect -1 -28 9 -24
rect 13 -28 23 -24
<< ntransistor >>
rect -5 -20 -3 -10
rect 5 -20 7 -10
rect 15 -20 17 -10
<< ptransistor >>
rect -5 8 -3 28
rect 5 8 7 28
rect 15 8 17 28
<< polycontact >>
rect -19 -2 -15 2
rect 0 1 4 5
rect 24 -2 28 2
<< ndcontact >>
rect -11 -14 -7 -10
rect -1 -20 3 -16
rect 9 -14 13 -10
rect 19 -20 23 -16
<< pdcontact >>
rect -11 8 -7 12
rect 19 24 23 28
<< psubstratepcontact >>
rect 9 -28 13 -24
<< nsubstratencontact >>
rect 3 34 7 38
<< labels >>
rlabel polycontact -19 -2 -15 2 7 vin_a
rlabel polycontact 0 1 4 5 7 vin_b
rlabel polycontact 24 -2 28 2 3 vin_c
rlabel metal1 -11 -8 -7 -4 7 vout
rlabel metal1 19 -28 23 -24 5 vss
rlabel metal1 17 34 21 38 1 vdd
<< end >>
